/* コア間割込み */

/* IPI を送出する */
[context("any")]
signature sIPISend{
    ER  sendIPI( [in]uint8_t ipino );
};

/* IPI を受信する */
[context("non-task"), callback]
signature sIPIMain{
    ER  main( void );
};

/*
 * コア間割込みを送る
 */
celltype tIPISenderUsingHSEM {
    /* User 側セルとの結合 */
    entry sIPISend          eIPISend;        /* コア間割込み発生させる */

    /* HSEM との結合 */
    call  sHSEM             cHSEM;          /* HSEM を使用して割込みを入れる */
    call  sHSEM             cHSEMGiantLock; /* HSEM を使用してGiantLock */

    attr {
        uint32_t           *ipi_bit_flag;   /* com_var.h の変数へのポインタ */
    };
};

/*
 * コア間割込みを受ける
 */
celltype tIPIReceiverUsingHSEM {
    /* User 側セルとの結合 */
    [optional]
        call  sIPIMain      cIPIMain[32];   /* コア間割込み受付ける */

    /* HSEM との結合 */
    call  sHSEM             cHSEMGiantLock; /* HSEM を使用してGiantLock */

    /* HSEM との結合 */
    entry siHSEMCallback    eCallback;      /* HSEM の割込みコールバック */

    attr {
        uint32_t           *ipi_bit_flag;   /* com_var.h の変数へのポインタ */
    };
};
