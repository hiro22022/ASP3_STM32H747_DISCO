/*
 *  TOPPERS/ASP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Advanced Standard Profile Kernel
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 *  Copyright (C) 2023 by hiro22022
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: target.cdl 648 2016-02-20 00:50:56Z ertl-honda $
 */
 
 import( "tIPI.cdl" );

 const uint32_t IPI_SysLog_4to7_NO  = 0;

/* Cortex M7 コアに割込みを送る */
[generate(CIfGenPlugin,"")]
cell tIPISenderUsingHSEM IPISender4to7 {
    /* HSEM との結合 */
    cHSEM = HSEMBody.eHSEM[HSEM_InterCoreInt_CM4_to_CM7];          /* HSEMBody.eHSEM[0] を使用 */
    cHSEMGiantLock = HSEMBody.eHSEM[HSEM_GiantLock];

    ipi_bit_flag = C_EXP( "&COM_IPI_4to7" );   /* com_var.h の変数へのポインタ */
};

/* Cortex M7 コアで割込みを受ける */
cell tIPIReceiverUsingHSEM IPIReceiver7to4 {
    /* HSEM との結合 */
    eCallback <= HSEMBody.cCallback[HSEM_InterCoreInt_CM7_to_CM4];	/* 逆結合 */
    cHSEMGiantLock = HSEMBody.eHSEM[HSEM_GiantLock];

    ipi_bit_flag = C_EXP( "&COM_IPI_7to4" );        /* com_var.h の変数へのポインタ */
};
