/*
 *		サンプルプログラム(1)のコンポーネント記述ファイル
 *
 *  $Id: sample1.cdl 839 2017-10-17 02:48:52Z ertl-hiro $
 */
/*
 *  カーネルオブジェクトの定義
 */
import(<kernel.cdl>);

/*
 *  ターゲット非依存のセルタイプの定義
 */
import("syssvc/tSerialPort.cdl");
import("syssvc/tSerialAdapter.cdl");
import("syssvc/tSysLog.cdl");
import("syssvc/tSysLogAdapter.cdl");
import("syssvc/tLogTask.cdl");
import("syssvc/tBanner.cdl");

/*
 *  ターゲット依存部の取り込み
 */
import("target.cdl");

/*
 *  「セルの組上げ記述」とは，"cell"で始まる行から，それに対応する"};"
 *  の行までのことを言う．
 */

/*
 *		システムログ機能のアダプタの組上げ記述
 *
 *  システムログ機能のアダプタは，C言語で記述されたコードから，TECSベー
 *  スのシステムログ機能を呼び出すためのセルである．システムログ機能の
 *  サービスコール（syslog，syslog_0〜syslog_5，t_perrorを含む）を呼び
 *  出さない場合には，以下のセルの組上げ記述を削除してよい．
 */
cell tSysLogAdapter SysLogAdapter {
	cSysLog = SysLog.eSysLog;
};

/*
 *		シリアルインタフェースドライバのアダプタの組上げ記述
 *
 *  シリアルインタフェースドライバのアダプタは，C言語で記述されたコー
 *  ドから，TECSベースのシリアルインタフェースドライバを呼び出すための
 *  セルである．シリアルインタフェースドライバのサービスコールを呼び出
 *  さない場合には，以下のセルの組上げ記述を削除してよい．
 */
cell tSerialAdapter SerialAdapter {
	cSerialPort[0] = SerialPort1.eSerialPort;
};

/*
 *		システムログ機能の組上げ記述
 *
 *  システムログ機能を外す場合には，以下のセルの組上げ記述を削除し，コ
 *  ンパイルオプションに-DTOPPERS_OMIT_SYSLOGを追加すればよい．ただし，
 *  システムログタスクはシステムログ機能を使用するため，それも外すこと
 *  が必要である．また，システムログ機能のアダプタも外さなければならな
 *  い．tecsgenが警告メッセージを出すが，無視してよい．
 */
cell tSysLog SysLog {
	logBufferSize = 32;					/* ログバッファのサイズ */
	initLogMask = C_EXP("LOG_UPTO(LOG_NOTICE)");
										/* ログバッファに記録すべき重要度 */
	initLowMask = C_EXP("LOG_UPTO(LOG_EMERG)");
									   	/* 低レベル出力すべき重要度 */
	/* 低レベル出力との結合 */
	cPutLog = PutLogTarget.ePutLog;
};

/*
 *		シリアルインタフェースドライバの組上げ記述
 *
 *  シリアルインタフェースドライバを外す場合には，以下のセルの組上げ記
 *  述を削除すればよい．ただし，システムログタスクはシリアルインタフェー
 *  スドライバを使用するため，それも外すことが必要である．また，シリア
 *  ルインタフェースドライバのアダプタも外さなければならない．
 */
cell tSerialPort SerialPort1 {
	receiveBufferSize = 256;			/* 受信バッファのサイズ */
	sendBufferSize    = 256;			/* 送信バッファのサイズ */

	/* ターゲット依存部との結合 */
	cSIOPort = SIOPortTarget1.eSIOPort;
	eiSIOCBR <= SIOPortTarget1.ciSIOCBR;	/* コールバック */
};

/*
 *		システムログタスクの組上げ記述
 *
 *  システムログタスクを外す場合には，以下のセルの組上げ記述を削除すれ
 *  ばよい．
 */
cell tLogTask LogTask {
	priority  = 3;					/* システムログタスクの優先度 */
	stackSize = LogTaskStackSize;	/* システムログタスクのスタックサイズ */

	/* シリアルインタフェースドライバとの結合 */
	cSerialPort        = SerialPort1.eSerialPort;
	cnSerialPortManage = SerialPort1.enSerialPortManage;

	/* システムログ機能との結合 */
	cSysLog = SysLog.eSysLog;

	/* 低レベル出力との結合 */
	cPutLog = PutLogTarget.ePutLog;
};

/*
 *		カーネル起動メッセージ出力の組上げ記述
 *
 *  カーネル起動メッセージの出力を外す場合には，以下のセルの組上げ記述
 *  を削除すればよい．
 */
cell tBanner Banner {
	/* 属性の設定 */
	targetName      = BannerTargetName;
	copyrightNotice = BannerCopyrightNotice;
};

/*
 * HSEM
 */
[singleton]
celltype tHSEM1Hanlder{
	entry siHSEMCallback eCallback;
	call  sHSEM    cHSEM;
};
cell tHSEM1Hanlder HSEM1Handler {
	eCallback <= HSEMBody.cCallback[0];	/* 逆結合 */
	cHSEM = HSEMBody.eHSEM[0];
};
